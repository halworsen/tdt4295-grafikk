// BRAM_SDP_MACRO: Simple Dual Port RAM
// 7 Series
// Xilinx HDL Libraries Guide, version 2012.2
///////////////////////////////////////////////////////////////////////
//  READ_WIDTH | BRAM_SIZE |  READ Depth | RDADDR Width |            //
// WRITE_WIDTH |           | WRITE Depth | WRADDR Width | WE Width   //
// ============|===========|=============|==============|============//
//    37-72    | "36Kb"    | 512         |  9-bit       | 8-bit      //
//    19-36    | "36Kb"    | 1024        | 10-bit       | 4-bit      //
//    19-36    | "18Kb"    | 512         |  9-bit       | 4-bit      //
//    10-18    | "36Kb"    | 2048        | 11-bit       | 2-bit      //
//    10-18    | "18Kb"    | 1024        | 10-bit       | 2-bit      //
//      5-9    | "36Kb"    | 4096        | 12-bit       | 1-bit      //
//      5-9    | "18Kb"    | 2048        | 11-bit       | 1-bit      //
//      3-4    | "36Kb"    | 8192        | 13-bit       | 1-bit      //
//      3-4    | "18Kb"    | 4096        | 12-bit       | 1-bit      //
//        2    | "36Kb"    | 16384       | 14-bit       | 1-bit      //
//        2    | "18Kb"    | 8192        | 13-bit       | 1-bit      //
//        1    | "36Kb"    | 32768       | 15-bit       | 1-bit      //
//        1    | "18Kb"    | 16384       | 14-bit       | 1-bit      //
///////////////////////////////////////////////////////////////////////

`default_nettype none
`timescale 1ns / 1ps

// BRAM_SDP_MACRO is documented in Xilinx UG472

module Bram #(
    // See table above fot the correct configuration
    parameter BRAM_SIZE="36Kb",   // BRAM size
    parameter WIDTH=1,
    //parameter DEPTH=2048,
    parameter DEPTH=32768,
    localparam ADDRW=$clog2(DEPTH),
    localparam INIT_FILE=""
) (
    input  wire logic clk_read,        // read clock
    input  wire logic clk_write,        // write clock
    input  wire logic reset,
    input  wire logic read_enable,
    input  wire logic write_enable,
    input  wire logic read_out_reg_en,
    input  wire logic writeport_enable,

    input  wire logic [ADDRW-1:0] read_addr,
    input  wire logic [ADDRW-1:0] write_addr,
    input  wire logic [WIDTH-1:0] data_in,        // data in
    output wire logic [WIDTH-1:0] data_out        // data out
    );

BRAM_SDP_MACRO #(
    .BRAM_SIZE(BRAM_SIZE), // Target BRAM, "18Kb" or "36Kb"
    .DEVICE("7SERIES"), // Target device: "7SERIES"
    .WRITE_WIDTH(WIDTH), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
    .READ_WIDTH(WIDTH), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
    .DO_REG(0), // Optional output register (0 or 1)
    .INIT_FILE(INIT_FILE),
    .SIM_COLLISION_CHECK("ALL"), // Collision check enable "ALL", "WARNING_ONLY",
    // "GENERATE_X_ONLY" or "NONE"
    .SRVAL(72'h00000000000000), // Set/Reset value forr port output
    .INIT(72'h08080808080808), // Initial values on output port
    .WRITE_MODE("WRITE_FIRST"), // Specify "READ_FIRST" forr same clock or synchronous clocks
    // Specify "WRITE_FIRST forr asynchronous clocks on ports
    //.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    // The next set of INIT_xx are valid when configured as 36Kb
    //.INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    //.INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    // The next set of INITP_xx are forr the parity bits
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    // The next set of INITP_xx are valid when configured as 36Kb
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_SDP_MACRO_inst (
    .DO(data_out),             // Output read data port, width defined by READ_WIDTH parameter
    .DI(data_in),             // Input write data port, width defined by WRITE_WIDTH parameter
    .RDADDR(read_addr),  // Input read address, width defined by read port depth
    .RDCLK(clk_read),    // 1-bit input read clock
    .RDEN(read_enable),  // 1-bit input read port enable
    .REGCE(read_out_reg_en),       // 1-bit input read output register enable
    .RST(reset),         // 1-bit input reset
    .WE(write_enable),   // Input write enable, width defined by write port depth
    .WRADDR(write_addr), // Input write address, width defined by write port depth
    .WRCLK(clk_write),   // 1-bit input write clock
    .WREN(writeport_enable)          // 1-bit input write port enable
);
// End of BRAM_SDP_MACRO_inst instantiation
endmodule
